`include "alu_interface.sv"


package pack;

	import p_headers::*;
	
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	
	`include "ALU_cfg.svh"
	`include "ALU_sequence_item.svh"
	`include "ALU_sequence.svh"
	`include "ALU_sequencer.svh"
	`include "ALU_driver.svh"
	`include "ALU_monitor.svh"
	`include "ALU_agent.svh"
	`include "ALU_scoreboard.svh"
	`include "ALU_coverage_collector.svh"
	`include "ALU_env.svh"
	`include "ALU_test.svh"
	
endpackage : pack


