/*######################################################################
## Class Name: Instruction_signed_min_sequence  
## Engineer : Omnia Mohamed
## Date: May 2025
## Description: 
    .This sequence is used to put min signed values in all registers using lui instruction. 
######################################################################*/
class Instruction_signed_min_sequence extends Instruction_base_Sequence;
    `uvm_object_utils(Instruction_signed_min_sequence)
    int num_transactions=31;
    Instruction_Seq_Item item;
    int count=0;
    function new(string name="Instruction_signed_min_sequence");
        super.new(name);
    endfunction
    virtual task body();
        super.body();
    endtask
    virtual task randomize_item();
        
        repeat(num_transactions)begin
            count=count+1;
            item=Instruction_Seq_Item::type_id::create("item");
            start_item(item);
            `uvm_info("Instruction_signed_min_sequence","seq is starting now",UVM_MEDIUM)
            
            assert(item.randomize() with{instruction_type==u_type;
					 utype==lui; imm==32'h8000_0000;
                                         rd==count;rs1==0;})
            else `uvm_fatal("Instruction_signed_min_sequence","Randomization Failed")
            `uvm_info("Instruction_signed_min_sequence","seq is randomized",UVM_MEDIUM)
            `uvm_info("Instruction_signed_min_sequence", item.sprint(),UVM_HIGH)
            `uvm_info("Instruction_signed_min_sequence","seq is finishing",UVM_MEDIUM)
            if(count==31)
                count=0;
            finish_item(item);
            
        end
    endtask
endclass
